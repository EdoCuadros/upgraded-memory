-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
-- Created on Sat Nov 05 12:25:22 2022

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SM2 IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        input2 : IN STD_LOGIC := '0';
        input3 : IN STD_LOGIC := '0';
        output1 : OUT STD_LOGIC
    );
END SM2;

ARCHITECTURE BEHAVIOR OF SM2 IS
    TYPE type_fstate IS (state1,state2,state3,state4,state5,state6,state7,state8);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,input2,input3)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            output1 <= '0';
        ELSE
            output1 <= '0';
            CASE fstate IS
                WHEN state1 =>
                    IF (((input2 = '1') AND (input3 = '0'))) THEN
                        reg_fstate <= state3;
                    ELSIF (((input2 = '1') AND (input3 = '1'))) THEN
                        reg_fstate <= state7;
                    ELSIF (((input2 = '0') AND (input3 = '0'))) THEN
                        reg_fstate <= state2;
                    ELSIF (((input2 = '0') AND (input3 = '1'))) THEN
                        reg_fstate <= state8;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;
                WHEN state2 =>
                    IF (((input2 = '0') AND (input3 = '0'))) THEN
                        reg_fstate <= state3;
                    ELSIF (((input2 = '1') AND (input3 = '0'))) THEN
                        reg_fstate <= state4;
                    ELSIF (((input2 = '0') AND (input3 = '1'))) THEN
                        reg_fstate <= state1;
                    ELSIF (((input2 = '1') AND (input3 = '1'))) THEN
                        reg_fstate <= state8;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    output1 <= '1';
                WHEN state3 =>
                    IF (((input2 = '0') AND (input3 = '0'))) THEN
                        reg_fstate <= state4;
                    ELSIF (((input2 = '0') AND (input3 = '1'))) THEN
                        reg_fstate <= state2;
                    ELSIF (((input2 = '1') AND (input3 = '0'))) THEN
                        reg_fstate <= state5;
                    ELSIF (((input2 = '1') AND (input3 = '1'))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;
                WHEN state4 =>
                    IF (((input2 = '1') AND (input3 = '0'))) THEN
                        reg_fstate <= state6;
                    ELSIF (((input2 = '0') AND (input3 = '1'))) THEN
                        reg_fstate <= state3;
                    ELSIF (((input2 = '0') AND (input3 = '0'))) THEN
                        reg_fstate <= state5;
                    ELSIF (((input2 = '1') AND (input3 = '1'))) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state4;
                    END IF;
                WHEN state5 =>
                    IF (((input2 = '0') AND (input3 = '0'))) THEN
                        reg_fstate <= state6;
                    ELSIF (((input2 = '1') AND (input3 = '0'))) THEN
                        reg_fstate <= state7;
                    ELSIF (((input2 = '0') AND (input3 = '1'))) THEN
                        reg_fstate <= state4;
                    ELSIF (((input2 = '1') AND (input3 = '1'))) THEN
                        reg_fstate <= state3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state5;
                    END IF;
                WHEN state6 =>
                    IF (((input2 = '0') AND (input3 = '0'))) THEN
                        reg_fstate <= state7;
                    ELSIF (((input2 = '1') AND (input3 = '1'))) THEN
                        reg_fstate <= state4;
                    ELSIF (((input2 = '0') AND (input3 = '1'))) THEN
                        reg_fstate <= state5;
                    ELSIF (((input2 = '1') AND (input3 = '0'))) THEN
                        reg_fstate <= state8;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state6;
                    END IF;
                WHEN state7 =>
                    IF (((input2 = '0') AND (input3 = '0'))) THEN
                        reg_fstate <= state8;
                    ELSIF (((input2 = '0') AND (input3 = '1'))) THEN
                        reg_fstate <= state6;
                    ELSIF (((input2 = '1') AND (input3 = '0'))) THEN
                        reg_fstate <= state1;
                    ELSIF (((input2 = '1') AND (input3 = '1'))) THEN
                        reg_fstate <= state5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state7;
                    END IF;
                WHEN state8 =>
                    IF (((input2 = '0') AND (input3 = '1'))) THEN
                        reg_fstate <= state7;
                    ELSIF (((input2 = '1') AND (input3 = '1'))) THEN
                        reg_fstate <= state6;
                    ELSIF (((input2 = '0') AND (input3 = '0'))) THEN
                        reg_fstate <= state1;
                    ELSIF (((input2 = '1') AND (input3 = '0'))) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state8;
                    END IF;
                WHEN OTHERS => 
                    output1 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
